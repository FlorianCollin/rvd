library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package my_cordic_rotati_pac is

  type vector_of_signed32 is ARRAY (NATURAL RANGE <>) OF signed(31 downto 0);

end package my_cordic_rotati_pac;

